module lab01_hello;
initial begin
	$display("Hello ModelSim!!");
end
endmodule